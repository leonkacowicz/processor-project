CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 20 30 90 10
176 80 1853 995
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
73 C:\Arquivos de programas\MicroCode Engineering\CircuitMaker 6 PRO\BOM.DAT
0 7
2 4 0.299301 0.500000
344 176 457 273
9508114 0
0
6 Title:
5 Name:
0
0
0
83
13 Logic Switch~
5 335 153 0 10 11
0 16 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-4 -16 10 -8
5 RESET
-14 -27 21 -19
0
0
25 *0=0V 1=5V

%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3765 0 0
2
42761.9 0
0
8 2-In OR~
219 1009 709 0 3 22
0 5 4 3
0
0 0 624 512
5 74F32
-18 -24 17 -16
4 U28C
-2 -25 26 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
3234 0 0
2
42761.9 1
0
10 2-In NAND~
219 1035 666 0 3 22
0 7 6 5
0
0 0 624 0
5 74F00
-10 -24 25 -16
4 U38C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 5 0
1 U
4155 0 0
2
42761.9 2
0
8 2-In OR~
219 966 639 0 3 22
0 9 8 6
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U28B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
6535 0 0
2
42761.9 3
0
9 2-In AND~
219 1039 630 0 3 22
0 6 7 10
0
0 0 624 692
5 74F08
-18 -24 17 -16
4 U34C
-17 -25 11 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 9 0
1 U
4527 0 0
2
42761.9 4
0
10 3-In NAND~
219 1559 365 0 4 22
0 49 11 50 51
0
0 0 624 512
5 74F10
-18 -28 17 -20
4 U42B
-11 -25 17 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 70
65 0 0 0 3 2 11 0
1 U
7899 0 0
2
42761.9 5
0
10 2-In NAND~
219 1424 353 0 3 22
0 109 108 9
0
0 0 624 0
5 74F00
-10 -24 25 -16
4 U38B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 5 0
1 U
4273 0 0
2
5.8939e-315 0
0
5 SCOPE
12 807 713 0 1 11
0 13
0
0 0 57584 0
5 RESET
-18 -4 17 4
3 U41
-11 -14 10 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
4787 0 0
2
42761.9 6
0
5 7474~
219 755 761 0 6 22
0 14 16 15 14 147 13
0
0 0 4720 0
5 74F74
4 -60 39 -52
4 U46A
23 -61 51 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
65 0 0 512 2 1 12 0
1 U
7655 0 0
2
42761.9 7
0
7 74LS244
143 1183 541 0 18 37
0 32 31 30 29 28 27 26 25 24
23 22 21 20 19 18 17 33 33
0
0 0 13040 0
6 74F244
-21 -60 21 -52
3 U45
-10 -61 11 -53
0
16 DVCC=20;DGND=10;
153 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %17i %18i]

+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %17o %18o %9o %10o %11o %12o %13o %14o %15o %16o] %M
0
12 type:digital
5 DIP20
37

0 8 6 4 2 11 13 15 17 12
14 16 18 9 7 5 3 1 19 8
6 4 2 11 13 15 17 12 14 16
18 9 7 5 3 1 19 0
65 0 0 0 1 1 0 0
1 U
8701 0 0
2
42761.9 8
0
6 PROM32
80 771 1112 0 14 29
0 34 35 36 37 38 39 8 12 148
149 150 151 152 153
0
0 0 4848 0
6 PROM32
-21 -19 21 -11
3 U44
-10 -61 11 -53
19 PROM_UC_BANK1_EXTRA
-69 -81 64 -73
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]

+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 2 3 4 5 6 7 9 10
11 12 13 14 15 1 2 3 4 5
6 7 9 10 11 12 13 14 15 0
65 0 0 512 1 0 0 0
1 U
5237 0 0
2
5.8939e-315 5.26354e-315
0
IAIAIAIAIAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
6 PROM32
80 533 1094 0 14 29
0 40 35 36 37 38 39 8 12 154
155 156 157 158 159
0
0 0 4336 0
6 PROM32
-21 -19 21 -11
3 U43
-10 -61 11 -53
19 PROM_UC_BANK0_EXTRA
-69 -81 64 -73
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]

+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 2 3 4 5 6 7 9 10
11 12 13 14 15 1 2 3 4 5
6 7 9 10 11 12 13 14 15 0
65 0 0 512 1 0 0 0
1 U
7721 0 0
2
5.8939e-315 5.30499e-315
0
IAIAIAIAIAIAIAIAIAIAIAAAIAIAIAIAMAIAIAIAIAIAIAIAIAIAIAIAIAIAIAIA
10 3-In NAND~
219 991 1046 0 4 22
0 68 11 67 41
0
0 0 624 0
5 74F10
-18 -28 17 -20
4 U42A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 70
65 0 0 0 3 1 11 0
1 U
9207 0 0
2
5.8939e-315 5.32571e-315
0
5 SCOPE
12 1036 1034 0 1 11
0 41
0
0 0 57584 0
4 CPIO
-14 -4 14 4
3 U41
-11 -14 10 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
9139 0 0
2
5.8939e-315 5.34643e-315
0
5 SCOPE
12 1031 1006 0 1 11
0 42
0
0 0 57584 0
4 CPSP
-14 -4 14 4
3 U41
-11 -14 10 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
9685 0 0
2
5.8939e-315 5.3568e-315
0
5 SCOPE
12 1031 975 0 1 11
0 43
0
0 0 57584 0
5 CPRES
-18 -4 17 4
3 U41
-11 -14 10 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
552 0 0
2
5.8939e-315 5.36716e-315
0
5 SCOPE
12 1031 946 0 1 11
0 44
0
0 0 57584 0
4 CPAC
-14 -4 14 4
3 U41
-11 -14 10 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
9878 0 0
2
5.8939e-315 5.37752e-315
0
5 SCOPE
12 1032 915 0 1 11
0 45
0
0 0 57584 0
4 CPIR
-14 -4 14 4
3 U41
-11 -14 10 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3800 0 0
2
5.8939e-315 5.38788e-315
0
5 SCOPE
12 1033 883 0 1 11
0 46
0
0 0 57584 0
4 cppc
-14 -4 14 4
3 U41
-11 -14 10 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
6962 0 0
2
5.8939e-315 5.39306e-315
0
5 SCOPE
12 1028 853 0 1 11
0 47
0
0 0 57584 0
5 cpmar
-18 -4 17 4
3 U41
-11 -14 10 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
5318 0 0
2
5.8939e-315 5.39824e-315
0
5 SCOPE
12 810 631 0 1 11
0 15
0
0 0 57584 0
2 CK
-8 -4 6 4
3 U41
-11 -14 10 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
9967 0 0
2
5.8939e-315 5.40342e-315
0
9 Inverter~
13 1607 356 0 2 22
0 48 49
0
0 0 624 180
6 74LS04
-21 -19 21 -11
4 U21F
-8 -20 20 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 2 0
1 U
963 0 0
2
42761.9 9
0
7 74LS244
143 1594 437 0 18 37
0 2 58 57 56 55 54 53 52 24
23 22 21 20 19 18 17 51 51
0
0 0 13040 0
6 74F244
-21 -60 21 -52
3 U40
-10 -61 11 -53
0
16 DVCC=20;DGND=10;
153 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %17i %18i]

+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %17o %18o %9o %10o %11o %12o %13o %14o %15o %16o] %M
0
12 type:digital
5 DIP20
37

0 8 6 4 2 11 13 15 17 12
14 16 18 9 7 5 3 1 19 8
6 4 2 11 13 15 17 12 14 16
18 9 7 5 3 1 19 0
65 0 0 0 1 1 0 0
1 U
4933 0 0
2
42761.9 10
0
9 Inverter~
13 940 1056 0 2 22
0 50 67
0
0 0 624 692
6 74LS04
-21 -19 21 -11
4 U21D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 2 0
1 U
323 0 0
2
42761.9 11
0
9 Inverter~
13 1552 326 0 2 22
0 11 69
0
0 0 624 692
6 74LS04
-21 -19 21 -11
4 U21C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 2 0
1 U
5628 0 0
2
42761.9 12
0
10 2-In NAND~
219 1610 317 0 3 22
0 71 69 70
0
0 0 624 0
5 74F00
-10 -24 25 -16
4 U38A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 62
65 0 0 0 4 1 5 0
1 U
9659 0 0
2
42761.9 13
0
6 74LS85
106 1586 248 0 14 29
0 66 65 64 63 14 14 14 14 74
73 72 160 11 161
0
0 0 13296 0
5 74F85
-18 -52 17 -44
3 U37
-11 -62 10 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]

+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 1 0 0 0
1 U
7883 0 0
2
42761.9 14
0
6 74LS85
106 1586 157 0 14 29
0 62 61 60 59 14 14 14 14 2
14 2 74 73 72
0
0 0 13296 0
5 74F85
-18 -52 17 -44
3 U36
-11 -62 10 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]

+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 18
65 0 0 0 1 0 0 0
1 U
358 0 0
2
42761.9 15
0
9 Inverter~
13 806 843 0 2 22
0 40 34
0
0 0 624 180
6 74LS04
-21 -19 21 -11
4 U21B
-8 -20 20 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
5235 0 0
2
5.8939e-315 5.4086e-315
0
6 PROM32
80 772 1000 0 14 29
0 34 35 36 37 38 39 83 33 82
81 80 48 50 7
0
0 0 4848 0
6 PROM32
-21 -19 21 -11
3 U35
-10 -61 11 -53
17 PROM_UC_BANK1_LOW
-62 -81 57 -73
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]

+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 2 3 4 5 6 7 9 10
11 12 13 14 15 1 2 3 4 5
6 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
7974 0 0
2
5.8939e-315 5.41378e-315
0
OPHPPLPLNJAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
6 PROM32
80 772 904 0 14 29
0 34 35 36 37 38 39 90 4 89
88 87 86 85 84
0
0 0 4848 0
6 PROM32
-21 -19 21 -11
3 U27
-10 -61 11 -53
18 PROM_UC_BANK1_HIGH
-66 -81 60 -73
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]

+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 2 3 4 5 6 7 9 10
11 12 13 14 15 1 2 3 4 5
6 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
4538 0 0
2
5.8939e-315 5.41896e-315
0
BCMDIDIDACAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
9 2-In AND~
219 991 987 0 3 22
0 87 68 43
0
0 0 624 692
5 74F08
-18 -24 17 -16
4 U34B
-17 -25 11 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 9 0
1 U
346 0 0
2
5.8939e-315 5.42414e-315
0
9 2-In AND~
219 991 1017 0 3 22
0 86 68 42
0
0 0 624 692
5 74F08
-18 -24 17 -16
4 U34A
-17 -25 11 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
3638 0 0
2
5.8939e-315 5.42933e-315
0
9 2-In AND~
219 991 926 0 3 22
0 89 68 45
0
0 0 624 692
5 74F08
-18 -24 17 -16
4 U33D
-17 -25 11 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 7 0
1 U
3628 0 0
2
5.8939e-315 5.43192e-315
0
9 2-In AND~
219 991 957 0 3 22
0 88 68 44
0
0 0 624 692
5 74F08
-18 -24 17 -16
4 U33C
-17 -25 11 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
5164 0 0
2
5.8939e-315 5.43451e-315
0
9 2-In AND~
219 991 896 0 3 22
0 3 68 46
0
0 0 624 692
5 74F08
-18 -24 17 -16
4 U33B
-17 -25 11 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
8570 0 0
2
5.8939e-315 5.4371e-315
0
9 2-In AND~
219 991 865 0 3 22
0 90 68 47
0
0 0 624 692
5 74F08
-18 -24 17 -16
4 U33A
-17 -25 11 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
8125 0 0
2
5.8939e-315 5.43969e-315
0
5 7474~
219 947 819 0 6 22
0 14 14 92 91 91 68
0
0 0 4720 0
5 74F74
4 -60 39 -52
4 U26B
23 -61 51 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 10 12 11 13 8 9 4 2 3
1 6 5 10 12 11 13 8 9 122
65 0 0 0 2 2 4 0
1 U
3154 0 0
2
5.8939e-315 0
0
6 PROM32
80 1387 494 0 14 29
0 2 2 32 31 30 29 162 163 94
95 96 97 98 99
0
0 0 4848 0
6 PROM32
-21 -19 21 -11
3 U32
-10 -61 11 -53
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]

+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 2 3 4 5 6 7 9 10
11 12 13 14 15 1 2 3 4 5
6 7 9 10 11 12 13 14 15 0
65 0 0 512 1 0 0 0
1 U
7583 0 0
2
5.8939e-315 5.26354e-315
0
CJAGBLBOBGAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
5 7425~
219 1352 344 0 6 22
0 107 106 105 104 14 109
0
0 0 624 0
4 7425
-14 -24 14 -16
4 U18A
-6 19 22 27
0
15 DVCC=14;DGND=7;
69 %D [%14bi %7bi %1i %2i %3i %4i %5i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 5 4 2 1 3 6 5 4 2
1 3 6 9 10 12 13 11 8 0
0 6 0
65 0 0 0 2 1 1 0
1 U
3912 0 0
2
5.8939e-315 5.30499e-315
0
5 7425~
219 1353 390 0 6 22
0 103 102 101 100 14 108
0
0 0 624 0
4 7425
-14 -24 14 -16
4 U18B
-6 19 22 27
0
15 DVCC=14;DGND=7;
69 %D [%14bi %7bi %1i %2i %3i %4i %5i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 9 10 12 13 11 8 5 4 2
1 3 6 9 10 12 13 11 8 0
0 6 0
65 0 0 0 2 2 1 0
1 U
8479 0 0
2
5.8939e-315 5.32571e-315
0
7 74LS181
132 1392 258 0 22 45
0 96 97 98 99 103 102 101 100 20
19 18 17 94 25 110 164 165 166 114
113 112 111
0
0 0 4848 0
6 74F181
-21 -69 21 -61
3 U17
-11 -70 10 -62
0
16 DVCC=24;DGND=12;
192 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i]

+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 3 4 5 6 19 21 23 2 18
20 22 1 7 8 16 14 17 15 13
11 10 9 3 4 5 6 19 21 23
2 18 20 22 1 7 8 16 14 17
15 13 11 10 9 0
65 0 0 512 1 0 0 0
1 U
3587 0 0
2
5.8939e-315 5.34643e-315
0
7 74LS181
132 1392 136 0 22 45
0 96 97 98 99 107 106 105 104 24
23 22 21 110 95 167 168 169 170 118
117 116 115
0
0 0 4848 0
6 74F181
-21 -69 21 -61
3 U15
-11 -70 10 -62
0
16 DVCC=24;DGND=12;
192 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i]

+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 3 4 5 6 19 21 23 2 18
20 22 1 7 8 16 14 17 15 13
11 10 9 3 4 5 6 19 21 23
2 18 20 22 1 7 8 16 14 17
15 13 11 10 9 0
65 0 0 512 1 0 0 0
1 U
5881 0 0
2
5.8939e-315 5.3568e-315
0
6 PROM32
80 539 88 0 14 29
0 119 63 62 61 60 59 24 23 22
21 20 19 18 17
0
0 0 4848 0
6 PROM32
-21 -19 21 -11
3 U31
-10 -61 11 -53
15 PROM_PROG_BANK0
-55 -81 50 -73
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]

+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 2 3 4 5 6 7 9 10
11 12 13 14 15 1 2 3 4 5
6 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
8486 0 0
2
42761.9 16
0
AFAEAEAAAAPPABGCACABABGBBKGCBIABADCKACGEAKGBBIABABGDAAGCBKGBAIAB
6 PROM32
80 539 184 0 14 29
0 120 63 62 61 60 59 24 23 22
21 20 19 18 17
0
0 0 4848 0
6 PROM32
-21 -19 21 -11
2 U2
-7 -61 7 -53
15 PROM_PROG_BANK1
-55 -81 50 -73
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]

+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 2 3 4 5 6 7 9 10
11 12 13 14 15 1 2 3 4 5
6 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
9939 0 0
2
42761.9 17
0
AMGDAAGBAIABABGBAEAMACABABGBBKGCBIABADEIACGEAKGBBIABABGDAHGDABPP
6 PROM32
80 539 280 0 14 29
0 121 63 62 61 60 59 24 23 22
21 20 19 18 17
0
0 0 4848 0
6 PROM32
-21 -19 21 -11
3 U29
-10 -61 11 -53
15 PROM_PROG_BANK2
-55 -81 50 -73
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]

+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 2 3 4 5 6 7 9 10
11 12 13 14 15 1 2 3 4 5
6 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
5351 0 0
2
42761.9 18
0
AAGBAIABABGBAECOAGAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAMM
7 74LS138
19 522 510 0 14 29
0 66 65 64 14 2 48 79 78 77
76 75 121 120 119
0
0 0 4848 0
6 74F138
-21 -61 21 -53
2 U6
-7 -71 7 -63
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]

+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 1 1 0 0
1 U
3216 0 0
2
42761.9 19
0
6 1K RAM
79 539 386 0 20 41
0 2 2 66 65 64 63 62 61 60
59 24 23 22 21 20 19 18 17 70
50
0
0 0 4848 0
5 RAM1K
-17 -19 18 -11
2 U1
-7 -70 7 -62
0
16 DVCC=22;DGND=11;
214 %D [%22bi %11bi  %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i %19i %20i]

+ [%22bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o  %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o] %M
0
12 type:digital
5 DIP22
41

0 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 0
65 0 0 0 1 0 0 0
1 U
7970 0 0
2
42761.9 20
0
10 8-In NAND~
219 590 487 0 9 19
0 14 14 14 79 78 77 76 75 71
0
0 0 624 0
5 74F30
-18 -24 17 -16
3 U19
-12 -44 9 -36
0
15 DVCC=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]

+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 1 2 3 4 5 6 11 12 8
1 2 3 4 5 6 11 12 8 0
65 0 0 0 1 0 0 0
1 U
7862 0 0
2
42761.9 21
0
12 Hex Display~
7 167 164 0 16 19
10 104 105 106 107 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 57184 0
4 1MEG
-15 -42 13 -34
3 ACh
-11 -38 10 -30
3 ACh
-10 -38 11 -30
0
50 %DA %1 0 %V

%DB %2 0 %V

%DC %3 0 %V

%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3440 0 0
2
42761.9 22
0
12 Hex Display~
7 199 164 0 18 19
10 100 101 102 103 0 0 0 0 0
0 1 1 1 1 1 1 1 8
0
0 0 55136 0
4 1MEG
-15 -42 13 -34
3 ACL
-11 -38 10 -30
3 ACL
-10 -39 11 -31
0
50 %DA %1 0 %V

%DB %2 0 %V

%DC %3 0 %V

%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
9128 0 0
2
42761.9 23
0
12 Hex Display~
7 119 165 0 18 19
10 137 136 135 134 0 0 0 0 0
0 1 1 1 1 1 1 1 8
0
0 0 54112 0
4 1MEG
-15 -42 13 -34
3 PCL
-11 -38 10 -30
3 PCL
-8 -38 13 -30
0
50 %DA %1 0 %V

%DB %2 0 %V

%DC %3 0 %V

%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3143 0 0
2
42761.9 24
0
12 Hex Display~
7 87 165 0 18 19
10 133 132 131 130 0 0 0 0 0
0 1 1 0 1 1 0 1 2
0
0 0 55136 0
4 1MEG
-15 -42 13 -34
3 PCh
-12 -38 9 -30
3 PCh
-10 -37 11 -29
0
50 %DA %1 0 %V

%DB %2 0 %V

%DC %3 0 %V

%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
374 0 0
2
42761.9 25
0
12 Hex Display~
7 162 276 0 18 19
10 63 64 65 66 0 0 0 0 0
0 1 0 1 1 1 1 1 6
0
0 0 55136 0
4 1MEG
-15 -42 13 -34
4 REGh
-14 -38 14 -30
4 REGh
-14 -37 14 -29
0
50 %DA %1 0 %V

%DB %2 0 %V

%DC %3 0 %V

%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3302 0 0
2
42761.9 26
0
12 Hex Display~
7 86 275 0 16 19
10 21 22 23 24 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 55136 0
4 1MEG
-15 -42 13 -34
5 busDh
-18 -38 17 -30
5 busDh
-20 -37 15 -29
0
50 %DA %1 0 %V

%DB %2 0 %V

%DC %3 0 %V

%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3949 0 0
2
42761.9 27
0
12 Hex Display~
7 118 275 0 18 19
10 17 18 19 20 0 0 0 0 0
0 1 1 1 1 1 1 1 8
0
0 0 55136 0
4 1MEG
-15 -42 13 -34
5 busDL
-18 -38 17 -30
5 busDL
-13 -36 22 -28
0
50 %DA %1 0 %V

%DB %2 0 %V

%DC %3 0 %V

%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
4216 0 0
2
42761.9 28
0
12 Hex Display~
7 198 276 0 18 19
10 59 60 61 62 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 55136 0
4 1MEG
-15 -42 13 -34
4 REGl
-15 -38 13 -30
4 REGl
-13 -38 15 -30
0
50 %DA %1 0 %V

%DB %2 0 %V

%DC %3 0 %V

%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
5936 0 0
2
42761.9 29
0
12 Hex Display~
7 86 384 0 16 19
10 29 30 31 32 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 55136 0
4 1MEG
-15 -42 13 -34
3 IRh
-11 -38 10 -30
3 IRh
-11 -39 10 -31
0
50 %DA %1 0 %V

%DB %2 0 %V

%DC %3 0 %V

%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
822 0 0
2
42761.9 30
0
12 Hex Display~
7 118 384 0 18 19
10 25 26 27 28 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 55136 0
4 1MEG
-15 -42 13 -34
3 IRL
-11 -38 10 -30
3 IRL
-10 -41 11 -33
0
50 %DA %1 0 %V

%DB %2 0 %V

%DC %3 0 %V

%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
6911 0 0
2
42761.9 31
0
12 Hex Display~
7 197 383 0 16 19
10 129 128 127 126 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 54112 0
4 1MEG
-15 -42 13 -34
3 SPL
-11 -38 10 -30
3 SPl
-10 -40 11 -32
0
50 %DA %1 0 %V

%DB %2 0 %V

%DC %3 0 %V

%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
674 0 0
2
42761.9 32
0
12 Hex Display~
7 165 383 0 16 19
10 125 124 123 122 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 55136 0
4 1MEG
-15 -42 13 -34
3 SPh
-11 -38 10 -30
3 SPh
-10 -39 11 -31
0
50 %DA %1 0 %V

%DB %2 0 %V

%DC %3 0 %V

%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3906 0 0
2
42761.9 33
0
14 Ascii Display~
172 136 592 0 42 44
0 23 22 21 20 19 18 17 41 0
0 8224 8224 8224 8224 8224 8224 8224 8224 8224
8224 8224 8224 8224 8224 8224 8224 8224 8224 8224
8224 8224 8224 8224 8224 8224 8224 8224 8224 8224
8224 8224 8224
0
0 0 21088 512
4 1MEG
-15 -42 13 -34
7 DISPLAY
-22 -48 27 -40
0
0
102 %DA %1 0 %V

%DB %2 0 %V

%DC %3 0 %V

%DD %4 0 %V

%DE %5 0 %V

%DF %6 0 %V

%DG %7 0 %V

%DH %8 0 %V
0
0
0
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
82 0 0 0 1 0 0 0
4 DISP
3411 0 0
2
42761.9 34
0
10 Ascii Key~
169 139 492 0 11 12
0 52 53 54 55 56 57 58 171 0
0 74
0
0 0 4656 0
0
7 Teclado
-24 -34 25 -26
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 512 1 0 0 0
3 KBD
4757 0 0
2
42761.9 35
0
7 74LS191
135 1187 218 0 14 29
0 2 42 13 12 14 14 14 2 145
172 126 127 128 129
0
0 0 4848 0
6 74F191
-21 -51 21 -43
3 U12
-11 -52 10 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]

+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 14 11 5 9 10 1 15 13
12 7 6 2 3 4 14 11 5 9
10 1 15 13 12 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
3199 0 0
2
42761.9 36
0
7 74LS191
135 1187 131 0 14 29
0 145 42 13 12 14 14 14 14 173
174 122 123 124 125
0
0 0 4848 0
6 74F191
-21 -51 21 -43
3 U22
-11 -52 10 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]

+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 14 11 5 9 10 1 15 13
12 7 6 2 3 4 14 11 5 9
10 1 15 13 12 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
8992 0 0
2
42761.9 37
0
7 74LS374
66 1187 440 0 34 37
0 118 117 116 115 114 113 112 111 24
23 22 21 20 19 18 17 81 43 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 1
0
0 0 13040 0
6 74F374
-21 -60 21 -52
3 U16
-11 -61 10 -53
0
16 DVCC=20;DGND=10;
153 %D [%20bi %10bi %17i %18i %1i %2i %3i %4i %5i %6i %7i %8i]

+ [%20bo %17o %18o %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o] %M
0
12 type:digital
5 DIP20
37

0 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 1 11 18
17 14 13 8 7 4 3 19 16 15
12 9 6 5 2 1 11 0
65 0 0 0 1 1 0 0
1 U
8789 0 0
2
42761.9 38
0
7 74LS374
66 750 162 0 37 37
0 24 23 22 21 20 19 18 17 66
65 64 63 62 61 60 59 2 47 0
0 0 0 0 0 0 0 0 0 0
0 1 1 0 0 0 0 1
0
0 0 13040 0
6 74F374
-21 -60 21 -52
2 U3
-7 -61 7 -53
0
16 DVCC=20;DGND=10;
153 %D [%20bi %10bi %17i %18i %1i %2i %3i %4i %5i %6i %7i %8i]

+ [%20bo %17o %18o %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o] %M
0
12 type:digital
5 DIP20
37

0 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 1 11 18
17 14 13 8 7 4 3 19 16 15
12 9 6 5 2 1 11 0
65 0 0 0 1 1 0 0
1 U
552 0 0
2
42761.9 39
0
7 74LS163
126 763 278 0 14 29
0 14 146 46 10 24 23 22 21 13
175 130 131 132 133
0
0 0 13040 0
7 74F163A
-25 -51 24 -43
2 U4
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]

+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 7 10 2 9 6 5 4 3 1
15 11 12 13 14 7 10 2 9 6
5 4 3 1 15 11 12 13 14 0
65 0 0 512 1 1 0 0
1 U
6515 0 0
2
42761.9 40
0
7 74LS163
126 763 370 0 14 29
0 14 14 46 10 20 19 18 17 13
146 134 135 136 137
0
0 0 13040 0
7 74F163A
-25 -51 24 -43
2 U5
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]

+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 7 10 2 9 6 5 4 3 1
15 11 12 13 14 7 10 2 9 6
5 4 3 1 15 11 12 13 14 0
65 0 0 0 1 1 0 0
1 U
3712 0 0
2
42761.9 41
0
7 74LS244
143 772 483 0 18 37
0 130 131 132 133 134 135 136 137 24
23 22 21 20 19 18 17 83 83
0
0 0 13040 0
6 74F244
-21 -60 21 -52
2 U7
-7 -61 7 -53
0
16 DVCC=20;DGND=10;
153 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %17i %18i]

+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %17o %18o %9o %10o %11o %12o %13o %14o %15o %16o] %M
0
12 type:digital
5 DIP20
37

0 8 6 4 2 11 13 15 17 12
14 16 18 9 7 5 3 1 19 8
6 4 2 11 13 15 17 12 14 16
18 9 7 5 3 1 19 0
65 0 0 0 1 1 0 0
1 U
8666 0 0
2
42761.9 42
0
7 74LS374
66 979 156 0 37 37
0 24 23 22 21 20 19 18 17 32
31 30 29 28 27 26 25 2 45 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 1
0
0 0 13040 0
6 74F374
-21 -60 21 -52
2 U8
-7 -61 7 -53
0
16 DVCC=20;DGND=10;
153 %D [%20bi %10bi %17i %18i %1i %2i %3i %4i %5i %6i %7i %8i]

+ [%20bo %17o %18o %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o] %M
0
12 type:digital
5 DIP20
37

0 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 1 11 18
17 14 13 8 7 4 3 19 16 15
12 9 6 5 2 1 11 0
65 0 0 0 1 1 0 0
1 U
3783 0 0
2
42761.9 43
0
6 PROM32
80 979 251 0 14 29
0 2 2 28 27 26 25 176 177 93
138 139 140 141 142
0
0 0 4848 0
6 PROM32
-21 -19 21 -11
2 U9
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]

+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 2 3 4 5 6 7 9 10
11 12 13 14 15 1 2 3 4 5
6 7 9 10 11 12 13 14 15 0
65 0 0 512 1 0 0 0
1 U
9918 0 0
2
42761.9 44
0
ACAFAIAKAMAOBDBGBKBKBNBNCBAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
7 74LS374
66 980 378 0 34 37
0 24 23 22 21 20 19 18 17 107
106 105 104 103 102 101 100 2 44 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 1
0
0 0 13040 0
6 74F374
-21 -60 21 -52
3 U10
-11 -61 10 -53
0
16 DVCC=20;DGND=10;
153 %D [%20bi %10bi %17i %18i %1i %2i %3i %4i %5i %6i %7i %8i]

+ [%20bo %17o %18o %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o] %M
0
12 type:digital
5 DIP20
37

0 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 1 11 18
17 14 13 8 7 4 3 19 16 15
12 9 6 5 2 1 11 0
65 0 0 0 1 1 0 0
1 U
3957 0 0
2
42761.9 45
0
7 74LS244
143 980 473 0 18 37
0 107 106 105 104 103 102 101 100 24
23 22 21 20 19 18 17 82 82
0
0 0 13040 0
6 74F244
-21 -60 21 -52
3 U11
-10 -61 11 -53
0
16 DVCC=20;DGND=10;
153 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %17i %18i]

+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %17o %18o %9o %10o %11o %12o %13o %14o %15o %16o] %M
0
12 type:digital
5 DIP20
37

0 8 6 4 2 11 13 15 17 12
14 16 18 9 7 5 3 1 19 8
6 4 2 11 13 15 17 12 14 16
18 9 7 5 3 1 19 0
65 0 0 0 1 1 0 0
1 U
8927 0 0
2
42761.9 46
0
7 74LS244
143 1188 314 0 18 37
0 122 123 124 125 126 127 128 129 24
23 22 21 20 19 18 17 80 80
0
0 0 13040 0
6 74F244
-21 -60 21 -52
3 U14
-10 -61 11 -53
0
16 DVCC=20;DGND=10;
153 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %17i %18i]

+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %17o %18o %9o %10o %11o %12o %13o %14o %15o %16o] %M
0
12 type:digital
5 DIP20
37

0 8 6 4 2 11 13 15 17 12
14 16 18 9 7 5 3 1 19 8
6 4 2 11 13 15 17 12 14 16
18 9 7 5 3 1 19 0
65 0 0 0 1 1 0 0
1 U
383 0 0
2
42761.9 47
0
7 Ground~
168 369 114 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8709 0 0
2
42761.9 48
0
2 +V
167 369 79 0 1 3
0 14
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3348 0 0
2
42761.9 49
0
7 74LS163
126 533 693 0 14 29
0 14 144 15 85 2 2 93 138 143
178 179 180 40 35
0
0 0 13040 0
7 74F163A
-25 -51 24 -43
3 U13
-10 -52 11 -44
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]

+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 7 10 2 9 6 5 4 3 1
15 11 12 13 14 7 10 2 9 6
5 4 3 1 15 11 12 13 14 0
65 0 0 512 1 1 0 0
1 U
8524 0 0
2
42761.9 50
0
7 74LS163
126 533 779 0 14 29
0 14 14 15 85 139 140 141 142 143
144 36 37 38 39
0
0 0 13040 0
7 74F163A
-25 -51 24 -43
3 U23
-10 -52 11 -44
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]

+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 7 10 2 9 6 5 4 3 1
15 11 12 13 14 7 10 2 9 6
5 4 3 1 15 11 12 13 14 0
65 0 0 0 1 1 0 0
1 U
8230 0 0
2
42761.9 51
0
6 PROM32
80 533 900 0 14 29
0 40 35 36 37 38 39 90 4 89
88 87 86 85 84
0
0 0 4848 0
6 PROM32
-21 -19 21 -11
3 U24
-11 -61 10 -53
18 PROM_UC_BANK0_HIGH
-66 -81 60 -73
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]

+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 2 3 4 5 6 7 9 10
11 12 13 14 15 1 2 3 4 5
6 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
4728 0 0
2
42761.9 52
0
MDCBMDIDBCMDIDACMDBCMDACMDACMDCDIHADACAHIDACMDIDIDBCMDALBCMDIDAL
6 PROM32
80 533 996 0 14 29
0 40 35 36 37 38 39 83 33 82
81 80 48 50 7
0
0 0 4336 0
6 PROM32
-21 -19 21 -11
3 U25
-10 -61 11 -53
17 PROM_UC_BANK0_LOW
-62 -81 57 -73
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]

+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 2 3 4 5 6 7 9 10
11 12 13 14 15 1 2 3 4 5
6 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
5697 0 0
2
42761.9 53
0
HPPLHPPLPLHPPLNJHPPLHPPLHPPKHPPLPHHJLOPPPHPKHPPLPLPLHPPLOPHPPLPL
9 2-In AND~
219 541 632 0 3 22
0 84 13 143
0
0 0 624 692
5 74F08
-18 -24 17 -16
4 U20B
-17 -25 11 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3849 0 0
2
42761.9 54
0
7 Pulser~
4 753 653 0 10 12
0 181 182 15 92 0 0 10 10 6
8
0
0 0 4656 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3356 0 0
2
42761.9 55
0
642
3 -867069182 3 0 0 4224 0 2 0 0 379 2
982 709
898 709
2 -13547956 4 0 0 4096 0 2 0 0 378 2
1028 718
1097 718
3 1 5 0 0 12416 0 3 2 0 0 4
1062 666
1066 666
1066 700
1028 700
2 0 6 0 0 8320 0 3 0 0 8 3
1011 675
1005 675
1005 639
1 0 7 0 0 4096 0 3 0 0 9 2
1011 657
1011 621
2 -13552231 8 0 0 4096 0 4 0 0 379 2
953 648
898 648
1 -29 9 0 0 4224 0 4 0 0 379 2
953 630
898 630
1 3 6 0 0 0 0 5 4 0 0 2
1015 639
999 639
2 -182887 7 0 0 4224 0 5 0 0 379 2
1015 621
898 621
3 -10173107 10 0 0 4096 0 5 0 0 378 2
1060 630
1097 630
2 -158568 11 0 0 4224 0 6 0 0 121 2
1585 365
1673 365
7 -13552231 8 0 0 4224 0 12 0 0 443 2
565 1067
647 1067
8 -9332851 12 0 0 4224 0 12 0 0 443 2
565 1076
647 1076
7 -13552231 8 0 0 0 0 11 0 0 398 2
803 1085
881 1085
8 -9332851 12 0 0 0 0 11 0 0 398 2
803 1094
881 1094
1 0 13 0 0 0 0 8 0 0 20 2
807 725
807 725
4 1 14 0 0 4096 0 9 0 0 399 2
755 773
673 773
1 1 14 0 0 0 0 9 0 0 399 2
755 698
673 698
3 -3303 15 0 0 4096 0 9 0 0 399 2
731 743
673 743
6 -616971363 13 0 0 4224 0 9 0 0 398 2
779 725
881 725
2 -149731 16 0 0 4096 0 9 0 0 399 2
731 725
673 725
-3264 16 17 0 0 12288 0 0 10 512 0 4
1267 585
1252 585
1252 586
1215 586
-3263 15 18 0 0 12288 0 0 10 512 0 4
1267 576
1252 576
1252 577
1215 577
-3262 14 19 0 0 12288 0 0 10 512 0 4
1267 567
1252 567
1252 568
1215 568
-3261 13 20 0 0 12288 0 0 10 512 0 4
1267 558
1252 558
1252 559
1215 559
-3260 12 21 0 0 12288 0 0 10 512 0 4
1267 540
1252 540
1252 541
1215 541
-3259 11 22 0 0 12288 0 0 10 512 0 4
1267 531
1252 531
1252 532
1215 532
-3258 10 23 0 0 12288 0 0 10 512 0 4
1267 522
1252 522
1252 523
1215 523
-3257 9 24 0 0 12288 0 0 10 512 0 4
1267 513
1252 513
1252 514
1215 514
8 -186688 25 0 0 4096 0 10 0 0 513 2
1151 586
1104 586
7 -186687 26 0 0 4096 0 10 0 0 513 2
1151 577
1104 577
6 -186686 27 0 0 4096 0 10 0 0 513 2
1151 568
1104 568
5 -186685 28 0 0 4096 0 10 0 0 513 2
1151 559
1104 559
4 -186684 29 0 0 4096 0 10 0 0 513 2
1151 541
1104 541
3 -186683 30 0 0 4096 0 10 0 0 513 2
1151 532
1104 532
2 -186682 31 0 0 4096 0 10 0 0 513 2
1151 523
1104 523
1 -186681 32 0 0 4096 0 10 0 0 513 2
1151 514
1104 514
18 -10427237 33 0 0 4096 0 10 0 0 513 2
1145 550
1104 550
17 -10427237 33 0 0 0 0 10 0 0 513 2
1145 505
1104 505
1 0 34 0 0 8192 0 11 0 0 149 3
733 1076
716 1076
716 964
2 -8863100 35 0 0 4096 0 11 0 0 399 2
739 1112
673 1112
3 -8863101 36 0 0 4096 0 11 0 0 399 2
739 1121
673 1121
4 -8863102 37 0 0 4096 0 11 0 0 399 2
739 1130
673 1130
5 -8863103 38 0 0 4096 0 11 0 0 399 2
739 1139
673 1139
6 -8863104 39 0 0 4096 0 11 0 0 399 2
739 1148
673 1148
2 -8863100 35 0 0 0 0 12 0 0 444 2
501 1094
436 1094
3 -8863101 36 0 0 0 0 12 0 0 444 2
501 1103
436 1103
4 -8863102 37 0 0 0 0 12 0 0 444 2
501 1112
436 1112
5 -8863103 38 0 0 0 0 12 0 0 444 2
501 1121
436 1121
6 -8863104 39 0 0 0 0 12 0 0 444 2
501 1130
436 1130
1 -8863099 40 0 0 4096 0 12 0 0 444 2
495 1058
436 1058
1 0 41 0 0 4096 0 14 0 0 107 2
1036 1046
1036 1055
1 0 42 0 0 4096 0 15 0 0 177 2
1031 1018
1031 1017
1 0 43 0 0 0 0 16 0 0 178 2
1031 987
1031 987
1 0 44 0 0 4096 0 17 0 0 179 2
1031 958
1031 957
1 0 45 0 0 4096 0 18 0 0 180 2
1032 927
1032 926
1 0 46 0 0 4096 0 19 0 0 181 2
1033 895
1033 896
1 0 47 0 0 0 0 20 0 0 182 2
1028 865
1028 865
1 0 15 0 0 0 0 21 0 0 397 2
810 643
810 644
1 -149731 16 0 0 4224 0 1 0 0 469 2
347 153
406 153
1 -864984170 48 0 0 4096 0 22 0 0 121 2
1628 356
1673 356
2 1 49 0 0 4224 0 22 6 0 0 2
1592 356
1585 356
3 -2336 50 0 0 4224 0 6 0 0 121 2
1585 374
1673 374
17 0 51 0 0 4096 0 23 0 0 65 2
1556 401
1534 401
4 18 51 0 0 4224 0 6 23 0 0 3
1534 365
1534 446
1556 446
9 -3257 24 0 0 4096 0 23 0 0 121 2
1626 410
1673 410
10 -3258 23 0 0 4096 0 23 0 0 121 2
1626 419
1673 419
11 -3259 22 0 0 4096 0 23 0 0 121 2
1626 428
1673 428
12 -3260 21 0 0 4096 0 23 0 0 121 2
1626 437
1673 437
13 -3261 20 0 0 4096 0 23 0 0 121 2
1626 455
1673 455
14 -3262 19 0 0 4096 0 23 0 0 121 2
1626 464
1673 464
15 -3263 18 0 0 4096 0 23 0 0 121 2
1626 473
1673 473
16 -3264 17 0 0 4096 0 23 0 0 121 2
1626 482
1673 482
8 -2944 52 0 0 4224 0 23 0 0 448 2
1562 482
1513 482
7 -2943 53 0 0 4224 0 23 0 0 448 2
1562 473
1513 473
6 -2942 54 0 0 4224 0 23 0 0 448 2
1562 464
1513 464
5 -2941 55 0 0 4224 0 23 0 0 448 2
1562 455
1513 455
4 -2940 56 0 0 4224 0 23 0 0 448 2
1562 437
1513 437
3 -2939 57 0 0 4224 0 23 0 0 448 2
1562 428
1513 428
2 -2938 58 0 0 4224 0 23 0 0 448 2
1562 419
1513 419
1 0 2 0 0 4096 0 23 0 0 448 2
1562 410
1513 410
1 -3456 59 0 0 4096 0 57 0 0 376 2
207 300
207 335
2 -3455 60 0 0 4096 0 57 0 0 376 2
201 300
201 335
3 -3454 61 0 0 4096 0 57 0 0 376 2
195 300
195 335
4 -3453 62 0 0 4096 0 57 0 0 376 2
189 300
189 335
1 -3452 63 0 0 4096 0 54 0 0 376 2
171 300
171 335
2 -3451 64 0 0 4096 0 54 0 0 376 2
165 300
165 335
3 -3450 65 0 0 4096 0 54 0 0 376 2
159 300
159 335
4 -3449 66 0 0 4096 0 54 0 0 376 2
153 300
153 335
1 -2944 52 0 0 0 0 63 0 0 97 2
160 516
160 533
2 -2943 53 0 0 0 0 63 0 0 97 2
154 516
154 533
3 -2942 54 0 0 0 0 63 0 0 97 2
148 516
148 533
4 -2941 55 0 0 0 0 63 0 0 97 2
142 516
142 533
5 -2940 56 0 0 0 0 63 0 0 97 2
136 516
136 533
6 -2939 57 0 0 0 0 63 0 0 97 2
130 516
130 533
7 -2938 58 0 0 0 0 63 0 0 97 2
124 516
124 533
-215140 0 1 0 0 4128 0 0 0 0 0 2
91 533
202 533
8 -13527912 41 0 0 4096 0 62 0 0 106 2
226 623
263 623
7 -3264 17 0 0 0 0 62 0 0 106 2
220 615
263 615
6 -3263 18 0 0 0 0 62 0 0 106 2
220 606
263 606
5 -3262 19 0 0 0 0 62 0 0 106 2
220 597
263 597
4 -3261 20 0 0 0 0 62 0 0 106 2
220 588
263 588
3 -3260 21 0 0 0 0 62 0 0 106 2
220 579
263 579
2 -3259 22 0 0 0 0 62 0 0 106 2
220 570
263 570
1 -3258 23 0 0 0 0 62 0 0 106 2
220 561
263 561
-215140 0 1 0 0 4128 0 0 0 0 0 2
263 517
263 648
4 -13527912 41 0 0 8320 0 13 0 0 378 5
1018 1046
1018 1055
1082 1055
1082 1047
1097 1047
1 -2336 50 0 0 0 0 24 0 0 379 2
925 1056
898 1056
2 3 67 0 0 4224 0 24 13 0 0 3
961 1056
967 1056
967 1055
2 -158568 11 0 0 0 0 13 0 0 379 4
967 1046
913 1046
913 1047
898 1047
1 0 68 0 0 8192 0 13 0 0 193 3
967 1037
953 1037
953 1008
1 -158568 11 0 0 0 0 25 0 0 448 2
1537 326
1513 326
2 2 69 0 0 4224 0 25 26 0 0 2
1573 326
1586 326
3 -864963946 70 0 0 4096 0 26 0 0 121 2
1637 317
1673 317
1 -150890 71 0 0 4224 0 26 0 0 448 2
1586 308
1513 308
9 -150890 71 0 0 0 0 49 0 0 641 2
617 487
647 487
13 -158568 11 0 0 0 0 27 0 0 121 2
1618 275
1673 275
11 0 2 0 0 4096 0 28 0 0 121 2
1618 148
1673 148
9 0 2 0 0 0 0 28 0 0 121 2
1618 130
1673 130
10 1 14 0 0 0 0 28 0 0 121 2
1618 139
1673 139
-215140 0 1 0 0 4128 0 0 0 0 0 2
1673 81
1673 562
8 1 14 0 0 0 0 27 0 0 448 2
1554 284
1513 284
7 1 14 0 0 0 0 27 0 0 448 2
1554 275
1513 275
6 1 14 0 0 0 0 27 0 0 448 2
1554 266
1513 266
5 1 14 0 0 0 0 27 0 0 448 2
1554 257
1513 257
8 1 14 0 0 0 0 28 0 0 448 2
1554 193
1513 193
7 1 14 0 0 0 0 28 0 0 448 2
1554 184
1513 184
6 1 14 0 0 0 0 28 0 0 448 2
1554 175
1513 175
5 1 14 0 0 0 0 28 0 0 448 2
1554 166
1513 166
4 -3452 63 0 0 4096 0 27 0 0 448 2
1554 248
1513 248
3 -3451 64 0 0 4096 0 27 0 0 448 2
1554 239
1513 239
2 -3450 65 0 0 4096 0 27 0 0 448 2
1554 230
1513 230
1 -3449 66 0 0 4096 0 27 0 0 448 2
1554 221
1513 221
4 -3456 59 0 0 4096 0 28 0 0 448 2
1554 157
1513 157
3 -3455 60 0 0 4096 0 28 0 0 448 2
1554 148
1513 148
2 -3454 61 0 0 4096 0 28 0 0 448 2
1554 139
1513 139
1 -3453 62 0 0 4096 0 28 0 0 448 2
1554 130
1513 130
14 11 72 0 0 8320 0 28 27 0 0 4
1618 193
1636 193
1636 239
1618 239
13 10 73 0 0 8320 0 28 27 0 0 4
1618 184
1631 184
1631 230
1618 230
12 9 74 0 0 8320 0 28 27 0 0 4
1618 175
1626 175
1626 221
1618 221
2 0 14 0 0 0 0 49 0 0 142 2
566 465
554 465
3 0 14 0 0 0 0 49 0 0 307 3
566 474
554 474
554 456
8 11 75 0 0 4224 0 49 47 0 0 2
566 519
560 519
7 10 76 0 0 4224 0 49 47 0 0 2
566 510
560 510
6 9 77 0 0 4224 0 49 47 0 0 2
566 501
560 501
5 8 78 0 0 4224 0 49 47 0 0 2
566 492
560 492
4 7 79 0 0 4224 0 49 47 0 0 2
566 483
560 483
1 0 34 0 0 0 0 31 0 0 149 2
734 868
716 868
2 1 34 0 0 8320 0 29 30 0 0 4
791 843
716 843
716 964
734 964
1 -8863099 40 0 0 0 0 29 0 0 398 2
827 843
881 843
14 -182887 7 0 0 0 0 30 0 0 398 2
804 1036
881 1036
13 -2336 50 0 0 0 0 30 0 0 398 2
804 1027
881 1027
12 -864984170 48 0 0 4096 0 30 0 0 398 2
804 1018
881 1018
11 -10426599 80 0 0 4096 0 30 0 0 398 2
804 1009
881 1009
10 -667307108 81 0 0 4096 0 30 0 0 398 2
804 1000
881 1000
9 -10427764 82 0 0 4096 0 30 0 0 398 2
804 991
881 991
8 -10427237 33 0 0 4096 0 30 0 0 398 2
804 982
881 982
7 -10426804 83 0 0 4096 0 30 0 0 398 2
804 973
881 973
14 -613296244 84 0 0 4096 0 31 0 0 398 2
804 940
881 940
13 -749103220 85 0 0 4096 0 31 0 0 398 2
804 931
881 931
12 -13547751 86 0 0 4096 0 31 0 0 398 2
804 922
881 922
11 -867060836 87 0 0 4096 0 31 0 0 398 2
804 913
881 913
10 -13548916 88 0 0 4096 0 31 0 0 398 2
804 904
881 904
9 -13548389 89 0 0 4096 0 31 0 0 398 2
804 895
881 895
8 -13547956 4 0 0 4096 0 31 0 0 398 2
804 886
881 886
7 -867081573 90 0 0 4096 0 31 0 0 398 2
804 877
881 877
2 -8863100 35 0 0 4096 0 30 0 0 399 2
740 1000
673 1000
3 -8863101 36 0 0 4096 0 30 0 0 399 2
740 1009
673 1009
4 -8863102 37 0 0 4096 0 30 0 0 399 2
740 1018
673 1018
5 -8863103 38 0 0 4096 0 30 0 0 399 2
740 1027
673 1027
6 -8863104 39 0 0 4096 0 30 0 0 399 2
740 1036
673 1036
2 -8863100 35 0 0 0 0 31 0 0 399 2
740 904
673 904
3 -8863101 36 0 0 0 0 31 0 0 399 2
740 913
673 913
4 -8863102 37 0 0 0 0 31 0 0 399 2
740 922
673 922
5 -8863103 38 0 0 0 0 31 0 0 399 2
740 931
673 931
6 -8863104 39 0 0 0 0 31 0 0 399 2
740 940
673 940
3 -13527271 42 0 0 4224 0 33 0 0 378 2
1012 1017
1097 1017
3 -865750116 43 0 0 4224 0 32 0 0 378 2
1012 987
1097 987
3 -13528436 44 0 0 4224 0 35 0 0 378 2
1012 957
1097 957
3 -13527909 45 0 0 4224 0 34 0 0 378 2
1012 926
1097 926
3 -13527476 46 0 0 4224 0 36 0 0 378 2
1012 896
1097 896
3 -865770853 47 0 0 4224 0 37 0 0 378 2
1012 865
1097 865
1 -13547751 86 0 0 0 0 33 0 0 379 2
967 1026
898 1026
1 -867060836 87 0 0 0 0 32 0 0 379 2
967 996
898 996
1 -13548916 88 0 0 0 0 35 0 0 379 2
967 966
898 966
1 -13548389 89 0 0 0 0 34 0 0 379 2
967 935
898 935
1 -867069182 3 0 0 0 0 36 0 0 379 2
967 905
898 905
1 -867081573 90 0 0 0 0 37 0 0 379 2
967 874
898 874
2 0 68 0 0 0 0 32 0 0 193 2
967 978
953 978
2 0 68 0 0 0 0 35 0 0 193 2
967 948
953 948
2 0 68 0 0 0 0 34 0 0 193 2
967 917
953 917
2 0 68 0 0 0 0 36 0 0 193 2
967 887
953 887
2 0 68 0 0 8320 0 33 0 0 194 3
967 1008
953 1008
953 856
2 -211382 68 0 0 0 0 37 0 0 379 2
967 856
898 856
6 -211382 68 0 0 0 0 38 0 0 378 2
971 783
1097 783
5 4 91 0 0 8320 0 38 38 0 0 5
977 801
981 801
981 839
947 839
947 831
1 1 14 0 0 0 0 38 0 0 379 2
947 756
898 756
3 -211374 92 0 0 4096 0 38 0 0 379 2
923 801
898 801
2 1 14 0 0 0 0 38 0 0 379 2
923 783
898 783
9 -11947195 93 0 0 4224 0 72 0 0 565 2
1011 242
1077 242
13 -8863099 40 0 0 4224 0 78 0 0 443 2
565 720
647 720
9 -3305 94 0 0 4224 0 39 0 0 470 2
1419 485
1487 485
10 -42 95 0 0 4224 0 39 0 0 470 2
1419 494
1487 494
11 -2301 96 0 0 4224 0 39 0 0 470 2
1419 503
1487 503
12 -2302 97 0 0 4224 0 39 0 0 470 2
1419 512
1487 512
13 -2303 98 0 0 4224 0 39 0 0 470 2
1419 521
1487 521
14 -2304 99 0 0 4224 0 39 0 0 470 2
1419 530
1487 530
2 0 2 0 0 4096 0 39 0 0 471 2
1355 494
1294 494
3 -186681 32 0 0 4096 0 39 0 0 471 2
1355 503
1294 503
4 -186682 31 0 0 4096 0 39 0 0 471 2
1355 512
1294 512
5 -186683 30 0 0 4096 0 39 0 0 471 2
1355 521
1294 521
6 -186684 29 0 0 4096 0 39 0 0 471 2
1355 530
1294 530
1 0 2 0 0 0 0 39 0 0 471 2
1349 458
1294 458
4 -2304 99 0 0 0 0 42 0 0 471 2
1360 240
1294 240
3 -2303 98 0 0 0 0 42 0 0 471 2
1360 231
1294 231
2 -2302 97 0 0 0 0 42 0 0 471 2
1360 222
1294 222
1 -2301 96 0 0 0 0 42 0 0 471 2
1360 213
1294 213
3 -29 9 0 0 0 0 7 0 0 470 2
1451 353
1487 353
4 -220416 100 0 0 4096 0 41 0 0 471 2
1336 404
1294 404
3 -220415 101 0 0 4096 0 41 0 0 471 2
1336 395
1294 395
2 -220414 102 0 0 4096 0 41 0 0 471 2
1336 386
1294 386
1 -220413 103 0 0 4096 0 41 0 0 471 4
1336 377
1309 377
1309 378
1294 378
4 -220412 104 0 0 4096 0 40 0 0 471 2
1335 358
1294 358
3 -220411 105 0 0 4096 0 40 0 0 471 2
1335 349
1294 349
2 -220410 106 0 0 4096 0 40 0 0 471 2
1335 340
1294 340
1 -220409 107 0 0 4096 0 40 0 0 471 2
1335 331
1294 331
5 1 14 0 0 0 0 41 0 0 471 2
1358 369
1294 369
5 1 14 0 0 0 0 40 0 0 471 2
1357 323
1294 323
2 6 108 0 0 8320 0 7 41 0 0 4
1400 362
1396 362
1396 390
1392 390
1 6 109 0 0 4224 0 7 40 0 0 2
1400 344
1391 344
13 -3305 94 0 0 0 0 42 0 0 470 2
1424 213
1487 213
15 13 110 0 0 8320 0 42 43 0 0 4
1424 249
1442 249
1442 91
1424 91
22 -14067840 111 0 0 4224 0 42 0 0 470 2
1430 312
1487 312
21 -14067839 112 0 0 4224 0 42 0 0 470 2
1430 303
1487 303
20 -14067838 113 0 0 4224 0 42 0 0 470 2
1430 294
1487 294
19 -14067837 114 0 0 4224 0 42 0 0 470 2
1430 285
1487 285
22 -14067836 115 0 0 4224 0 43 0 0 470 2
1430 190
1487 190
21 -14067835 116 0 0 4224 0 43 0 0 470 2
1430 181
1487 181
20 -14067834 117 0 0 4224 0 43 0 0 470 2
1430 172
1487 172
19 -14067833 118 0 0 4224 0 43 0 0 470 2
1430 163
1487 163
12 -3264 17 0 0 4096 0 42 0 0 471 2
1354 312
1294 312
11 -3263 18 0 0 4096 0 42 0 0 471 2
1354 303
1294 303
10 -3262 19 0 0 4096 0 42 0 0 471 2
1354 294
1294 294
9 -3261 20 0 0 4096 0 42 0 0 471 2
1354 285
1294 285
12 -3260 21 0 0 4096 0 43 0 0 471 2
1354 190
1294 190
11 -3259 22 0 0 4096 0 43 0 0 471 2
1354 181
1294 181
10 -3258 23 0 0 4096 0 43 0 0 471 2
1354 172
1294 172
9 -3257 24 0 0 4096 0 43 0 0 471 2
1354 163
1294 163
8 -220416 100 0 0 4096 0 42 0 0 471 2
1354 276
1294 276
7 -220415 101 0 0 4096 0 42 0 0 471 2
1354 267
1294 267
6 -220414 102 0 0 4096 0 42 0 0 471 2
1354 258
1294 258
5 -220413 103 0 0 4096 0 42 0 0 471 2
1354 249
1294 249
8 -220412 104 0 0 4096 0 43 0 0 471 2
1354 154
1294 154
7 -220411 105 0 0 4096 0 43 0 0 471 2
1354 145
1294 145
6 -220410 106 0 0 4096 0 43 0 0 471 2
1354 136
1294 136
5 -220409 107 0 0 4096 0 43 0 0 471 2
1354 127
1294 127
14 -186688 25 0 0 4096 0 42 0 0 470 2
1424 222
1487 222
14 -42 95 0 0 0 0 43 0 0 470 2
1424 100
1487 100
4 -2304 99 0 0 0 0 43 0 0 471 2
1360 118
1294 118
3 -2303 98 0 0 0 0 43 0 0 471 2
1360 109
1294 109
2 -2302 97 0 0 0 0 43 0 0 471 2
1360 100
1294 100
1 -2301 96 0 0 0 0 43 0 0 471 2
1360 91
1294 91
1 -9599616 119 0 0 8192 0 44 0 0 642 3
501 52
501 79
438 79
7 -3257 24 0 0 4224 0 44 0 0 641 2
571 61
647 61
8 -3258 23 0 0 4224 0 44 0 0 641 2
571 70
647 70
9 -3259 22 0 0 4224 0 44 0 0 641 2
571 79
647 79
10 -3260 21 0 0 4224 0 44 0 0 641 2
571 88
647 88
11 -3261 20 0 0 4224 0 44 0 0 641 2
571 97
647 97
12 -3262 19 0 0 4224 0 44 0 0 641 2
571 106
647 106
13 -3263 18 0 0 4224 0 44 0 0 641 2
571 115
647 115
14 -3264 17 0 0 4224 0 44 0 0 641 2
571 124
647 124
2 -3452 63 0 0 4096 0 44 0 0 642 2
507 88
438 88
3 -3453 62 0 0 4096 0 44 0 0 642 2
507 97
438 97
4 -3454 61 0 0 4096 0 44 0 0 642 2
507 106
438 106
5 -3455 60 0 0 4096 0 44 0 0 642 2
507 115
438 115
6 -3456 59 0 0 4096 0 44 0 0 642 2
507 124
438 124
1 -9599615 120 0 0 4096 0 45 0 0 642 2
501 148
438 148
7 -3257 24 0 0 0 0 45 0 0 641 2
571 157
647 157
8 -3258 23 0 0 0 0 45 0 0 641 2
571 166
647 166
9 -3259 22 0 0 0 0 45 0 0 641 2
571 175
647 175
10 -3260 21 0 0 0 0 45 0 0 641 2
571 184
647 184
11 -3261 20 0 0 0 0 45 0 0 641 2
571 193
647 193
12 -3262 19 0 0 0 0 45 0 0 641 2
571 202
647 202
13 -3263 18 0 0 0 0 45 0 0 641 2
571 211
647 211
14 -3264 17 0 0 0 0 45 0 0 641 2
571 220
647 220
2 -3452 63 0 0 0 0 45 0 0 642 2
507 184
438 184
3 -3453 62 0 0 0 0 45 0 0 642 2
507 193
438 193
4 -3454 61 0 0 0 0 45 0 0 642 2
507 202
438 202
5 -3455 60 0 0 0 0 45 0 0 642 2
507 211
438 211
6 -3456 59 0 0 0 0 45 0 0 642 2
507 220
438 220
1 -9599614 121 0 0 4096 0 46 0 0 642 2
501 244
438 244
7 -3257 24 0 0 0 0 46 0 0 641 2
571 253
647 253
8 -3258 23 0 0 0 0 46 0 0 641 2
571 262
647 262
9 -3259 22 0 0 0 0 46 0 0 641 2
571 271
647 271
10 -3260 21 0 0 0 0 46 0 0 641 2
571 280
647 280
11 -3261 20 0 0 0 0 46 0 0 641 2
571 289
647 289
12 -3262 19 0 0 0 0 46 0 0 641 2
571 298
647 298
13 -3263 18 0 0 0 0 46 0 0 641 2
571 307
647 307
14 -3264 17 0 0 0 0 46 0 0 641 2
571 316
647 316
2 -3452 63 0 0 0 0 46 0 0 642 2
507 280
438 280
3 -3453 62 0 0 0 0 46 0 0 642 2
507 289
438 289
4 -3454 61 0 0 0 0 46 0 0 642 2
507 298
438 298
5 -3455 60 0 0 0 0 46 0 0 642 2
507 307
438 307
6 -3456 59 0 0 0 0 46 0 0 642 2
507 316
438 316
12 -9599614 121 0 0 4224 0 47 0 0 641 2
560 528
647 528
13 -9599615 120 0 0 4224 0 47 0 0 641 2
560 537
647 537
1 1 14 0 0 4224 0 49 0 0 642 2
566 456
438 456
6 -864984170 48 0 0 0 0 47 0 0 642 2
484 546
438 546
14 -9599616 119 0 0 4224 0 47 0 0 641 2
560 546
647 546
4 1 14 0 0 0 0 47 0 0 642 2
490 528
438 528
1 -3449 66 0 0 4096 0 47 0 0 642 2
490 483
438 483
2 -3450 65 0 0 4096 0 47 0 0 642 2
490 492
438 492
3 -3451 64 0 0 4096 0 47 0 0 642 2
490 501
438 501
0 5 2 0 0 0 0 0 47 642 0 2
438 537
484 537
20 -2336 50 0 0 0 0 48 0 0 641 2
577 359
647 359
19 -864963946 70 0 0 4224 0 48 0 0 641 2
577 350
647 350
11 -3257 24 0 0 0 0 48 0 0 641 2
571 368
647 368
12 -3258 23 0 0 0 0 48 0 0 641 2
571 377
647 377
13 -3259 22 0 0 0 0 48 0 0 641 2
571 386
647 386
14 -3260 21 0 0 0 0 48 0 0 641 2
571 395
647 395
15 -3261 20 0 0 0 0 48 0 0 641 2
571 404
647 404
16 -3262 19 0 0 0 0 48 0 0 641 2
571 413
647 413
17 -3263 18 0 0 0 0 48 0 0 641 2
571 422
647 422
18 -3264 17 0 0 0 0 48 0 0 641 2
571 431
647 431
2 0 2 0 0 4224 0 48 0 0 642 2
507 359
438 359
1 0 2 0 0 0 0 48 0 0 642 2
507 350
438 350
3 -3449 66 0 0 4096 0 48 0 0 642 2
507 368
438 368
4 -3450 65 0 0 4096 0 48 0 0 642 2
507 377
438 377
5 -3451 64 0 0 4096 0 48 0 0 642 2
507 386
438 386
6 -3452 63 0 0 0 0 48 0 0 642 2
507 395
438 395
7 -3453 62 0 0 0 0 48 0 0 642 2
507 404
438 404
8 -3454 61 0 0 0 0 48 0 0 642 2
507 413
438 413
9 -3455 60 0 0 0 0 48 0 0 642 2
507 422
438 422
10 -3456 59 0 0 0 0 48 0 0 642 2
507 431
438 431
4 -145849 122 0 0 4096 0 61 0 0 375 2
156 407
156 440
3 -145850 123 0 0 4096 0 61 0 0 375 2
162 407
162 440
2 -145851 124 0 0 4096 0 61 0 0 375 2
168 407
168 440
1 -145852 125 0 0 4096 0 61 0 0 375 2
174 407
174 440
4 -145853 126 0 0 4096 0 60 0 0 375 2
188 407
188 440
3 -145854 127 0 0 4096 0 60 0 0 375 2
194 407
194 440
2 -145855 128 0 0 4096 0 60 0 0 375 2
200 407
200 440
1 -145856 129 0 0 4096 0 60 0 0 375 2
206 407
206 440
4 -186681 32 0 0 0 0 58 0 0 375 2
77 408
77 440
3 -186682 31 0 0 0 0 58 0 0 375 2
83 408
83 440
2 -186683 30 0 0 0 0 58 0 0 375 2
89 408
89 440
1 -186684 29 0 0 0 0 58 0 0 375 2
95 408
95 440
4 -186685 28 0 0 0 0 59 0 0 375 2
109 408
109 440
3 -186686 27 0 0 0 0 59 0 0 375 2
115 408
115 440
2 -186687 26 0 0 0 0 59 0 0 375 2
121 408
121 440
1 -186688 25 0 0 0 0 59 0 0 375 2
127 408
127 440
4 -3257 24 0 0 0 0 55 0 0 376 2
77 299
77 335
3 -3258 23 0 0 0 0 55 0 0 376 2
83 299
83 335
2 -3259 22 0 0 0 0 55 0 0 376 2
89 299
89 335
1 -3260 21 0 0 0 0 55 0 0 376 2
95 299
95 335
4 -3261 20 0 0 0 0 56 0 0 376 2
109 299
109 335
3 -3262 19 0 0 0 0 56 0 0 376 2
115 299
115 335
2 -3263 18 0 0 0 0 56 0 0 376 2
121 299
121 335
1 -3264 17 0 0 0 0 56 0 0 376 2
127 299
127 335
4 -220409 107 0 0 0 0 50 0 0 377 2
158 188
158 228
3 -220410 106 0 0 0 0 50 0 0 377 2
164 188
164 228
2 -220411 105 0 0 0 0 50 0 0 377 2
170 188
170 228
1 -220412 104 0 0 0 0 50 0 0 377 2
176 188
176 228
4 -220413 103 0 0 0 0 51 0 0 377 2
190 188
190 228
3 -220414 102 0 0 0 0 51 0 0 377 2
196 188
196 228
2 -220415 101 0 0 0 0 51 0 0 377 2
202 188
202 228
1 -220416 100 0 0 0 0 51 0 0 377 2
208 188
208 228
4 -158969 130 0 0 4096 0 53 0 0 377 2
78 189
78 228
3 -158970 131 0 0 4096 0 53 0 0 377 2
84 189
84 228
2 -158971 132 0 0 4096 0 53 0 0 377 2
90 189
90 228
1 -158972 133 0 0 4096 0 53 0 0 377 2
96 189
96 228
4 -158973 134 0 0 4096 0 52 0 0 377 2
110 189
110 228
3 -158974 135 0 0 4096 0 52 0 0 377 2
116 189
116 228
2 -158975 136 0 0 4096 0 52 0 0 377 2
122 189
122 228
1 -158976 137 0 0 4096 0 52 0 0 377 2
128 189
128 228
-215140 0 1 0 0 32 0 0 0 0 0 2
242 440
59 440
-215140 0 1 0 0 32 0 0 0 0 0 2
240 335
59 335
-215140 0 1 0 0 32 0 0 0 0 0 2
240 228
57 228
-215140 0 1 0 0 4128 0 0 0 0 0 2
1097 602
1097 1089
-215140 0 1 0 0 32 0 0 0 0 0 2
898 607
898 1094
14 -182887 7 0 0 0 0 81 0 0 443 2
565 1032
647 1032
13 -2336 50 0 0 0 0 81 0 0 443 2
565 1023
647 1023
12 -864984170 48 0 0 4224 0 81 0 0 443 2
565 1014
647 1014
11 -10426599 80 0 0 4224 0 81 0 0 443 2
565 1005
647 1005
10 -667307108 81 0 0 4224 0 81 0 0 443 2
565 996
647 996
9 -10427764 82 0 0 4224 0 81 0 0 443 2
565 987
647 987
8 -10427237 33 0 0 4224 0 81 0 0 443 2
565 978
647 978
7 -10426804 83 0 0 4224 0 81 0 0 443 2
565 969
647 969
14 -613296244 84 0 0 4224 0 80 0 0 443 2
565 936
647 936
13 -749103220 85 0 0 4224 0 80 0 0 443 2
565 927
647 927
12 -13547751 86 0 0 4224 0 80 0 0 443 2
565 918
647 918
11 -867060836 87 0 0 4224 0 80 0 0 443 2
565 909
647 909
10 -13548916 88 0 0 4224 0 80 0 0 443 2
565 900
647 900
9 -13548389 89 0 0 4224 0 80 0 0 443 2
565 891
647 891
8 -13547956 4 0 0 4224 0 80 0 0 443 2
565 882
647 882
7 -867081573 90 0 0 4224 0 80 0 0 443 2
565 873
647 873
4 -211374 92 0 0 4224 0 83 0 0 398 2
783 653
881 653
3 -3303 15 0 0 4224 0 83 0 0 398 2
777 644
881 644
-215140 0 1 0 0 4128 0 0 0 0 0 2
881 607
881 1161
-215140 0 1 0 0 4256 0 0 0 0 0 2
673 601
673 1162
3 -3303 15 0 0 0 0 79 0 0 444 2
501 770
436 770
3 -3303 15 0 0 0 0 78 0 0 444 2
501 684
436 684
7 -11947195 93 0 0 0 0 78 0 0 444 2
501 720
436 720
6 0 2 0 0 0 0 78 0 0 444 2
501 711
436 711
5 0 2 0 0 0 0 78 0 0 444 2
501 702
436 702
8 -11947196 138 0 0 4096 0 78 0 0 444 2
501 729
436 729
5 -11947197 139 0 0 4096 0 79 0 0 444 2
501 788
436 788
6 -11947198 140 0 0 4096 0 79 0 0 444 2
501 797
436 797
7 -11947199 141 0 0 4096 0 79 0 0 444 2
501 806
436 806
8 -11947200 142 0 0 4096 0 79 0 0 444 2
501 815
436 815
10 -11947196 138 0 0 4224 0 72 0 0 565 2
1011 251
1077 251
11 -11947197 139 0 0 4224 0 72 0 0 565 2
1011 260
1077 260
12 -11947198 140 0 0 4224 0 72 0 0 565 2
1011 269
1077 269
13 -11947199 141 0 0 4224 0 72 0 0 565 2
1011 278
1077 278
14 -11947200 142 0 0 4224 0 72 0 0 565 2
1011 287
1077 287
2 -8863100 35 0 0 0 0 81 0 0 444 2
501 996
436 996
3 -8863101 36 0 0 0 0 81 0 0 444 2
501 1005
436 1005
4 -8863102 37 0 0 0 0 81 0 0 444 2
501 1014
436 1014
5 -8863103 38 0 0 0 0 81 0 0 444 2
501 1023
436 1023
6 -8863104 39 0 0 0 0 81 0 0 444 2
501 1032
436 1032
2 -8863100 35 0 0 0 0 80 0 0 444 2
501 900
436 900
3 -8863101 36 0 0 0 0 80 0 0 444 2
501 909
436 909
4 -8863102 37 0 0 0 0 80 0 0 444 2
501 918
436 918
5 -8863103 38 0 0 0 0 80 0 0 444 2
501 927
436 927
6 -8863104 39 0 0 0 0 80 0 0 444 2
501 936
436 936
1 -8863099 40 0 0 0 0 81 0 0 444 2
495 960
436 960
1 -8863099 40 0 0 0 0 80 0 0 444 2
495 864
436 864
9 0 143 0 0 4096 0 78 0 0 428 2
571 666
586 666
9 3 143 0 0 8320 0 79 82 0 0 4
571 752
586 752
586 632
562 632
1 -613296244 84 0 0 0 0 82 0 0 444 2
517 641
436 641
2 -616971363 13 0 0 0 0 82 0 0 444 2
517 623
436 623
14 -8863100 35 0 0 4224 0 78 0 0 443 2
565 729
647 729
11 -8863101 36 0 0 4224 0 79 0 0 443 2
565 788
647 788
12 -8863102 37 0 0 4224 0 79 0 0 443 2
565 797
647 797
13 -8863103 38 0 0 4224 0 79 0 0 443 2
565 806
647 806
14 -8863104 39 0 0 4224 0 79 0 0 443 2
565 815
647 815
2 1 14 0 0 0 0 79 0 0 444 2
501 761
436 761
4 -749103220 85 0 0 0 0 79 0 0 444 2
495 779
436 779
4 -749103220 85 0 0 0 0 78 0 0 444 2
495 693
436 693
2 -584005822 144 0 0 4096 0 78 0 0 444 2
501 675
436 675
10 -584005822 144 0 0 4224 0 79 0 0 443 2
565 779
647 779
1 1 14 0 0 0 0 78 0 0 444 2
501 666
436 666
1 1 14 0 0 0 0 79 0 0 444 2
501 752
436 752
-215140 0 1 0 0 32 0 0 0 0 0 2
647 601
647 1162
-215140 0 1 0 0 32 0 0 0 0 0 2
436 607
436 1161
1 0 2 0 0 0 0 64 0 0 513 2
1149 191
1104 191
1 -9648359 145 0 0 4224 0 65 0 0 513 2
1149 104
1104 104
2 -13527271 42 0 0 0 0 65 0 0 513 2
1155 113
1104 113
-215140 0 1 0 0 32 0 0 0 0 0 2
1513 82
1513 563
8 -14067840 111 0 0 0 0 66 0 0 513 2
1155 476
1104 476
7 -14067839 112 0 0 0 0 66 0 0 513 2
1155 467
1104 467
6 -14067838 113 0 0 0 0 66 0 0 513 2
1155 458
1104 458
5 -14067837 114 0 0 0 0 66 0 0 513 2
1155 449
1104 449
4 -14067836 115 0 0 0 0 66 0 0 513 2
1155 440
1104 440
3 -14067835 116 0 0 0 0 66 0 0 513 2
1155 431
1104 431
2 -14067834 117 0 0 0 0 66 0 0 513 2
1155 422
1104 422
1 -14067833 118 0 0 0 0 66 0 0 513 2
1155 413
1104 413
9 -3257 24 0 0 0 0 66 0 0 512 2
1219 413
1267 413
10 -3258 23 0 0 0 0 66 0 0 512 2
1219 422
1267 422
11 -3259 22 0 0 0 0 66 0 0 512 2
1219 431
1267 431
12 -3260 21 0 0 0 0 66 0 0 512 2
1219 440
1267 440
13 -3261 20 0 0 0 0 66 0 0 512 2
1219 449
1267 449
14 -3262 19 0 0 0 0 66 0 0 512 2
1219 458
1267 458
15 -3263 18 0 0 0 0 66 0 0 512 2
1219 467
1267 467
16 -3264 17 0 0 0 0 66 0 0 512 2
1219 476
1267 476
18 -865750116 43 0 0 0 0 66 0 0 512 2
1219 404
1267 404
17 -667307108 81 0 0 0 0 66 0 0 513 2
1149 404
1104 404
1 0 2 0 0 0 0 76 0 0 469 2
369 108
406 108
1 1 14 0 0 0 0 77 0 0 469 2
369 88
406 88
-215140 0 1 0 0 32 0 0 0 0 0 2
406 65
406 169
-215140 0 1 0 0 32 0 0 0 0 0 2
1487 81
1487 562
-215140 0 1 0 0 32 0 0 0 0 0 2
1294 78
1294 559
9 -3257 24 0 0 0 0 75 0 0 512 2
1220 287
1267 287
10 -3258 23 0 0 0 0 75 0 0 512 2
1220 296
1267 296
11 -3259 22 0 0 0 0 75 0 0 512 2
1220 305
1267 305
12 -3260 21 0 0 0 0 75 0 0 512 2
1220 314
1267 314
13 -3261 20 0 0 0 0 75 0 0 512 2
1220 332
1267 332
14 -3262 19 0 0 0 0 75 0 0 512 2
1220 341
1267 341
15 -3263 18 0 0 0 0 75 0 0 512 2
1220 350
1267 350
16 -3264 17 0 0 0 0 75 0 0 512 2
1220 359
1267 359
17 -10426599 80 0 0 0 0 75 0 0 513 2
1150 278
1104 278
18 -10426599 80 0 0 0 0 75 0 0 513 2
1150 323
1104 323
1 -145849 122 0 0 4224 0 75 0 0 513 2
1156 287
1104 287
2 -145850 123 0 0 4224 0 75 0 0 513 2
1156 296
1104 296
3 -145851 124 0 0 4224 0 75 0 0 513 2
1156 305
1104 305
4 -145852 125 0 0 4224 0 75 0 0 513 2
1156 314
1104 314
5 -145853 126 0 0 4224 0 75 0 0 513 2
1156 332
1104 332
6 -145854 127 0 0 4224 0 75 0 0 513 2
1156 341
1104 341
7 -145855 128 0 0 4224 0 75 0 0 513 2
1156 350
1104 350
8 -145856 129 0 0 4224 0 75 0 0 513 2
1156 359
1104 359
11 -145849 122 0 0 0 0 65 0 0 512 2
1219 140
1267 140
12 -145850 123 0 0 0 0 65 0 0 512 2
1219 149
1267 149
13 -145851 124 0 0 0 0 65 0 0 512 2
1219 158
1267 158
14 -145852 125 0 0 0 0 65 0 0 512 2
1219 167
1267 167
9 -9648359 145 0 0 0 0 64 0 0 512 2
1225 209
1267 209
11 -145853 126 0 0 0 0 64 0 0 512 2
1219 227
1267 227
12 -145854 127 0 0 0 0 64 0 0 512 2
1219 236
1267 236
13 -145855 128 0 0 0 0 64 0 0 512 2
1219 245
1267 245
14 -145856 129 0 0 0 0 64 0 0 512 2
1219 254
1267 254
3 -616971363 13 0 0 0 0 64 0 0 513 2
1149 209
1104 209
8 0 2 0 0 0 0 64 0 0 513 2
1155 254
1104 254
7 1 14 0 0 0 0 64 0 0 513 2
1155 245
1104 245
6 1 14 0 0 0 0 64 0 0 513 2
1155 236
1104 236
5 1 14 0 0 0 0 64 0 0 513 2
1155 227
1104 227
4 -9332851 12 0 0 0 0 64 0 0 513 2
1155 218
1104 218
2 -13527271 42 0 0 0 0 64 0 0 513 2
1155 200
1104 200
3 -616971363 13 0 0 0 0 65 0 0 513 2
1149 122
1104 122
8 1 14 0 0 0 0 65 0 0 513 2
1155 167
1104 167
7 1 14 0 0 0 0 65 0 0 513 2
1155 158
1104 158
6 1 14 0 0 0 0 65 0 0 513 2
1155 149
1104 149
5 1 14 0 0 0 0 65 0 0 513 2
1155 140
1104 140
4 -9332851 12 0 0 0 0 65 0 0 513 2
1155 131
1104 131
-215140 0 1 0 0 32 0 0 0 0 0 2
1267 78
1267 599
-215140 0 1 0 0 32 0 0 0 0 0 2
1104 77
1104 599
8 -220416 100 0 0 0 0 74 0 0 575 2
948 518
892 518
7 -220415 101 0 0 0 0 74 0 0 575 2
948 509
892 509
6 -220414 102 0 0 0 0 74 0 0 575 2
948 500
892 500
5 -220413 103 0 0 0 0 74 0 0 575 2
948 491
892 491
4 -220412 104 0 0 0 0 74 0 0 575 2
948 473
892 473
3 -220411 105 0 0 0 0 74 0 0 575 2
948 464
892 464
2 -220410 106 0 0 0 0 74 0 0 575 2
948 455
892 455
1 -220409 107 0 0 0 0 74 0 0 575 2
948 446
892 446
-3264 16 17 0 0 0 0 0 74 565 0 2
1077 518
1012 518
-3263 15 18 0 0 0 0 0 74 565 0 2
1077 509
1012 509
-3262 14 19 0 0 0 0 0 74 565 0 2
1077 500
1012 500
-3261 13 20 0 0 0 0 0 74 565 0 2
1077 491
1012 491
-3260 12 21 0 0 0 0 0 74 565 0 2
1077 473
1012 473
-3259 11 22 0 0 0 0 0 74 565 0 2
1077 464
1012 464
-3258 10 23 0 0 0 0 0 74 565 0 2
1077 455
1012 455
-3257 9 24 0 0 0 0 0 74 565 0 2
1077 446
1012 446
18 -10427764 82 0 0 0 0 74 0 0 575 2
942 482
892 482
17 -10427764 82 0 0 0 0 74 0 0 575 2
942 437
892 437
18 -13528436 44 0 0 0 0 73 0 0 565 2
1012 342
1077 342
17 0 2 0 0 0 0 73 0 0 575 2
942 342
892 342
1 -3257 24 0 0 0 0 73 0 0 575 2
948 351
892 351
2 -3258 23 0 0 0 0 73 0 0 575 2
948 360
892 360
3 -3259 22 0 0 0 0 73 0 0 575 2
948 369
892 369
4 -3260 21 0 0 0 0 73 0 0 575 2
948 378
892 378
5 -3261 20 0 0 0 0 73 0 0 575 2
948 387
892 387
6 -3262 19 0 0 0 0 73 0 0 575 2
948 396
892 396
7 -3263 18 0 0 0 0 73 0 0 575 2
948 405
892 405
8 -3264 17 0 0 0 0 73 0 0 575 2
948 414
892 414
9 -220409 107 0 0 4224 0 73 0 0 565 2
1012 351
1077 351
10 -220410 106 0 0 4224 0 73 0 0 565 2
1012 360
1077 360
11 -220411 105 0 0 4224 0 73 0 0 565 2
1012 369
1077 369
12 -220412 104 0 0 4224 0 73 0 0 565 2
1012 378
1077 378
13 -220413 103 0 0 4224 0 73 0 0 565 2
1012 387
1077 387
14 -220414 102 0 0 4224 0 73 0 0 565 2
1012 396
1077 396
15 -220415 101 0 0 4224 0 73 0 0 565 2
1012 405
1077 405
16 -220416 100 0 0 4224 0 73 0 0 565 2
1012 414
1077 414
3 -186685 28 0 0 4096 0 72 0 0 575 2
947 260
892 260
4 -186686 27 0 0 4096 0 72 0 0 575 2
947 269
892 269
5 -186687 26 0 0 4096 0 72 0 0 575 2
947 278
892 278
6 -186688 25 0 0 0 0 72 0 0 575 2
947 287
892 287
1 0 2 0 0 0 0 72 0 0 575 2
941 215
892 215
2 0 2 0 0 0 0 72 0 0 575 2
947 251
892 251
9 -186681 32 0 0 4224 0 71 0 0 565 2
1011 129
1077 129
10 -186682 31 0 0 4224 0 71 0 0 565 2
1011 138
1077 138
11 -186683 30 0 0 4224 0 71 0 0 565 2
1011 147
1077 147
12 -186684 29 0 0 4224 0 71 0 0 565 2
1011 156
1077 156
13 -186685 28 0 0 4224 0 71 0 0 565 2
1011 165
1077 165
14 -186686 27 0 0 4224 0 71 0 0 565 2
1011 174
1077 174
15 -186687 26 0 0 4224 0 71 0 0 565 2
1011 183
1077 183
16 -186688 25 0 0 4224 0 71 0 0 565 2
1011 192
1077 192
18 -13527909 45 0 0 0 0 71 0 0 565 2
1011 120
1077 120
-215140 0 1 0 0 32 0 0 0 0 0 2
1077 77
1077 558
1 -3257 24 0 0 0 0 71 0 0 575 2
947 129
892 129
2 -3258 23 0 0 0 0 71 0 0 575 2
947 138
892 138
3 -3259 22 0 0 0 0 71 0 0 575 2
947 147
892 147
4 -3260 21 0 0 0 0 71 0 0 575 2
947 156
892 156
5 -3261 20 0 0 0 0 71 0 0 575 2
947 165
892 165
6 -3262 19 0 0 0 0 71 0 0 575 2
947 174
892 174
7 -3263 18 0 0 0 0 71 0 0 575 2
947 183
892 183
8 -3264 17 0 0 0 0 71 0 0 575 2
947 192
892 192
17 0 2 0 0 0 0 71 0 0 575 2
941 120
892 120
-215140 0 1 0 0 32 0 0 0 0 0 2
892 73
892 554
-3260 12 21 0 0 0 0 0 70 630 0 2
867 483
804 483
-3259 11 22 0 0 0 0 0 70 630 0 2
867 474
804 474
-3258 10 23 0 0 0 0 0 70 630 0 2
867 465
804 465
-3257 9 24 0 0 0 0 0 70 630 0 2
867 456
804 456
-3264 16 17 0 0 0 0 0 70 630 0 2
867 528
804 528
-3263 15 18 0 0 0 0 0 70 630 0 2
867 519
804 519
-3262 14 19 0 0 0 0 0 70 630 0 2
867 510
804 510
-3261 13 20 0 0 0 0 0 70 630 0 2
867 501
804 501
18 -10426804 83 0 0 0 0 70 0 0 640 2
734 492
673 492
17 -10426804 83 0 0 0 0 70 0 0 640 2
734 447
673 447
1 -158969 130 0 0 4096 0 70 0 0 640 2
740 456
673 456
2 -158970 131 0 0 4096 0 70 0 0 640 2
740 465
673 465
3 -158971 132 0 0 4096 0 70 0 0 640 2
740 474
673 474
4 -158972 133 0 0 4096 0 70 0 0 640 2
740 483
673 483
5 -158973 134 0 0 4096 0 70 0 0 640 2
740 501
673 501
6 -158974 135 0 0 4096 0 70 0 0 640 2
740 510
673 510
7 -158975 136 0 0 4096 0 70 0 0 640 2
740 519
673 519
8 -158976 137 0 0 4096 0 70 0 0 640 2
740 528
673 528
11 -158973 134 0 0 4224 0 69 0 0 630 2
795 379
867 379
12 -158974 135 0 0 4224 0 69 0 0 630 2
795 388
867 388
13 -158975 136 0 0 4224 0 69 0 0 630 2
795 397
867 397
14 -158976 137 0 0 4224 0 69 0 0 630 2
795 406
867 406
8 -3264 17 0 0 0 0 69 0 0 640 2
731 406
673 406
7 -3263 18 0 0 0 0 69 0 0 640 2
731 397
673 397
6 -3262 19 0 0 0 0 69 0 0 640 2
731 388
673 388
5 -3261 20 0 0 0 0 69 0 0 640 2
731 379
673 379
4 -10173107 10 0 0 4224 0 69 0 0 640 2
725 370
673 370
9 -616971363 13 0 0 0 0 69 0 0 630 2
801 343
867 343
2 1 14 0 0 0 0 69 0 0 640 2
731 352
673 352
1 1 14 0 0 0 0 69 0 0 640 2
731 343
673 343
3 -13527476 46 0 0 0 0 69 0 0 640 2
731 361
673 361
10 -584006755 146 0 0 4224 0 69 0 0 630 2
795 370
867 370
11 -158969 130 0 0 4224 0 68 0 0 630 2
795 287
867 287
12 -158970 131 0 0 4224 0 68 0 0 630 2
795 296
867 296
13 -158971 132 0 0 4224 0 68 0 0 630 2
795 305
867 305
14 -158972 133 0 0 4224 0 68 0 0 630 2
795 314
867 314
5 -3257 24 0 0 0 0 68 0 0 640 2
731 287
673 287
6 -3258 23 0 0 0 0 68 0 0 640 2
731 296
673 296
7 -3259 22 0 0 0 0 68 0 0 640 2
731 305
673 305
8 -3260 21 0 0 0 0 68 0 0 640 2
731 314
673 314
4 -10173107 10 0 0 0 0 68 0 0 640 2
725 278
673 278
9 -616971363 13 0 0 0 0 68 0 0 630 2
801 251
867 251
3 -13527476 46 0 0 0 0 68 0 0 640 2
731 269
673 269
2 -584006755 146 0 0 0 0 68 0 0 640 2
731 260
673 260
1 1 14 0 0 0 0 68 0 0 640 2
731 251
673 251
16 -3456 59 0 0 4224 0 67 0 0 630 2
782 198
867 198
15 -3455 60 0 0 4224 0 67 0 0 630 2
782 189
867 189
14 -3454 61 0 0 4224 0 67 0 0 630 2
782 180
867 180
13 -3453 62 0 0 4224 0 67 0 0 630 2
782 171
867 171
12 -3452 63 0 0 4224 0 67 0 0 630 2
782 162
867 162
11 -3451 64 0 0 4224 0 67 0 0 630 2
782 153
867 153
10 -3450 65 0 0 4224 0 67 0 0 630 2
782 144
867 144
9 -3449 66 0 0 4224 0 67 0 0 630 2
782 135
867 135
18 -865770853 47 0 0 0 0 67 0 0 630 2
782 126
867 126
-215140 0 1 0 0 32 0 0 0 0 0 2
867 73
867 554
1 -3257 24 0 0 0 0 67 0 0 640 2
718 135
673 135
2 -3258 23 0 0 0 0 67 0 0 640 2
718 144
673 144
3 -3259 22 0 0 0 0 67 0 0 640 2
718 153
673 153
4 -3260 21 0 0 0 0 67 0 0 640 2
718 162
673 162
5 -3261 20 0 0 0 0 67 0 0 640 2
718 171
673 171
6 -3262 19 0 0 0 0 67 0 0 640 2
718 180
673 180
7 -3263 18 0 0 0 0 67 0 0 640 2
718 189
673 189
8 -3264 17 0 0 0 0 67 0 0 640 2
718 198
673 198
17 0 2 0 0 0 0 67 0 0 640 2
712 126
673 126
-215140 0 1 0 0 32 0 0 0 0 0 2
673 71
673 552
-215140 0 1 0 0 32 0 0 0 0 0 2
647 27
647 569
-215140 0 1 0 0 32 0 0 0 0 0 2
438 65
438 563
11
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 86
334 212 424 334
337 215 420 313
86 DECODIFICADOR 

DO BANCO DE 

MEMORIA:

0 -> ROM0

1 -> ROM1

2 -> ROM2

OUTROS -> RAM
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 19
405 580 541 599
409 583 536 596
19 UNIDADE DE CONTROLE
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 10
422 21 496 40
425 25 492 38
10 COMPUTADOR
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 3
738 96 763 114
740 98 760 110
3 MAR
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
743 222 761 240
745 224 758 236
2 PC
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
963 86 982 105
966 89 978 102
2 IR
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
969 310 989 329
972 313 985 326
2 AC
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
1172 64 1192 83
1175 68 1188 81
2 SP
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 3
1173 368 1200 387
1176 372 1196 385
3 RES
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 3
1379 54 1406 73
1382 57 1402 70
3 ALU
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 23
1310 418 1470 437
1313 421 1466 434
23 DECOD. DE FUNCAO DA ALU
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 1e-06 1e-07 1e-07
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
